-------------------------------------------------------------------------------
--
-- Title       : \EX- project\
-- Design      : b
-- Author      : Aubai
-- Company     : non
--
-------------------------------------------------------------------------------
--
-- File        : C:/Users/Aubai/Desktop/Digital Logic/VHDL - examlpes/EX- project.vhd
-- Generated   : Fri Jan  1 16:51:24 2021
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {\EX- project\} architecture {\EX- project\}}



entity \EX- project\ is
end \EX- project\;

--}} End of automatically maintained section

architecture \EX- project\ of \EX- project\ is
begin

	 -- enter your statements here --

end \EX- project\;
