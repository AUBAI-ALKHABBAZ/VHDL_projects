SIGNAL x : BIT ;
x <= '0' ;
SIGNAL y : BIT_VECTOR( 3 DOWNTO 0 ) ;
y <= "0111" ;

 SIGNAL w ; BIT_VECTOR ( 7 DOWNTO 0 ) ;
 w <= "0111010" ;
 
 