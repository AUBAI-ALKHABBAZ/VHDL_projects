SIGNAL a : STD_LOGIC ;
a <= "101111" ; -- decimal 47
a <= 0"57" ;   -- بل أوكتال
a <= x"2f"; -- ستاعشري
VARIABLE b : INTEGER ;
b <= 1300 ;
